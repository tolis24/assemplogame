library ieee;
use ieee.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity icon_rom is
port (countV : in std_logic_vector(9 downto 0);
		pointer : in std_logic_vector(3 downto 0);
		dataOut : out std_logic_vector(79 downto 0));
end icon_rom;

architecture RTL of icon_rom is

signal row : std_logic_vector(9 downto 0);
signal address : std_logic_vector(9 downto 0);

begin

process (countV)
begin 
	if unsigned(countV) < 60 then 
		row <= countV;
	elsif unsigned(countV) < 120 then
		row <= unsigned(countV) - 60;
	elsif unsigned(countV) < 180 then
		row <= unsigned(countV) - 120;
	elsif unsigned(countV) < 240 then
		row <= unsigned(countV) - 180;
	elsif unsigned(countV) < 300 then
		row <= unsigned(countV) - 240;
	elsif unsigned(countV) < 360 then
		row <= unsigned(countV) - 300;
	elsif unsigned(countV) < 420 then
		row <= unsigned(countV) - 360;
	elsif unsigned(countV) < 480 then
		row <= unsigned(countV) - 420;
	else
		row <= (others => '0');
	end if;
end process;

		
address(9 downto 6) <= pointer;
address(5 downto 0) <= row(5 downto 0);

process(address)
begin
case address is
-- 0
when "0000000000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000000001"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000000010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000000011"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000000100"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000000101"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000000110"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000000111"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000001000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000001001"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000001010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000001011"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000001100"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000001101"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000001110"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000001111"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000010000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000010001"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000010010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000010011"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000010100"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000010101"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000010110"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000010111"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000011000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000011001"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000011010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000011011"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000011100"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000011101"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000011110"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000011111"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000100000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000100001"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000100010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000100011"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000100100"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000100101"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000100110"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000100111"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000101000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000101001"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000101010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000101011"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000101100"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000101101"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000101110"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000101111"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000110000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000110001"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000110010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000110011"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000110100"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000110101"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000110110"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000110111"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000111000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000111001"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000111010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000111011"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";

--1
when "0001000000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0001000001"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0001000010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0001000011"=> dataOut <= "00000000000000000000000000000000000000001100000000000000000000000000000000000000";
when "0001000100"=> dataOut <= "00000000000000000000000000000000000000011110000000000000000000000000000000000000";
when "0001000101"=> dataOut <= "00000000000000000000000000000000000000111111000000000000000000000000000000000000";
when "0001000110"=> dataOut <= "00000000000000000000000000000000000001110011100000000000000000000000000000000000";
when "0001000111"=> dataOut <= "00000000000000000000000000000000000011100011100000000000000000000000000000000000";
when "0001001000"=> dataOut <= "00000000000000000000000000000000000111000001110000000000000000000000000000000000";
when "0001001001"=> dataOut <= "00000000000000000000000000000000001110000000111000000000000000000000000000000000";
when "0001001010"=> dataOut <= "00000000000000000000000000000000011100000000011100000000000000000000000000000000";
when "0001001011"=> dataOut <= "00000000000000000000000000000000111000000000001110000000000000000000000000000000";
when "0001001100"=> dataOut <= "00000000000000000000000000000001110000000000000111000000000000000000000000000000";
when "0001001101"=> dataOut <= "00000000000000000000000000000011100000000000000011100000000000000000000000000000";
when "0001001110"=> dataOut <= "00000000000000000000000000000111000000000000000001110000000000000000000000000000";
when "0001001111"=> dataOut <= "00000000000000000000000000001110000000000000000000111000000000000000000000000000";
when "0001010000"=> dataOut <= "00000000000000000000000000011100000000000000000000011100000000000000000000000000";
when "0001010001"=> dataOut <= "00000000000000000000000000111000000000000000000000001110000000000000000000000000";
when "0001010010"=> dataOut <= "00000000000000000000000001110000000000000000000000000111000000000000000000000000";
when "0001010011"=> dataOut <= "00000000000000000000000011100000000000000000000000000011100000000000000000000000";
when "0001010100"=> dataOut <= "00000000000000000000000111000000000000000000000000000001110000000000000000000000";
when "0001010101"=> dataOut <= "00000000000000000000001110000000000000000000000000000000111000000000000000000000";
when "0001010110"=> dataOut <= "00000000000000000000011100000000000000000000000000000000011100000000000000000000";
when "0001010111"=> dataOut <= "00000000000000000000111000000000000000000000000000000000001110000000000000000000";
when "0001011000"=> dataOut <= "00000000000000000001110000000000000000000000000000000000000111000000000000000000";
when "0001011001"=> dataOut <= "00000000000000000011100000000000000000000000000000000000000011100000000000000000";
when "0001011010"=> dataOut <= "00000000000000000111000000000000000000000000000000000000000001110000000000000000";
when "0001011011"=> dataOut <= "00000000000000001110000000000000000000000000000000000000000000111000000000000000";
when "0001011100"=> dataOut <= "00000000000000011100000000000000000000000000000000000000000000011100000000000000";
when "0001011101"=> dataOut <= "00000000000000111000000000000000000000000000000000000000000000001110000000000000";
when "0001011110"=> dataOut <= "00000000000001110000000000000000000000000000000000000000000000000111000000000000"; --center
when "0001011111"=> dataOut <= "00000000000000111000000000000000000000000000000000000000000000001110000000000000";
when "0001100000"=> dataOut <= "00000000000000011100000000000000000000000000000000000000000000011100000000000000";
when "0001100001"=> dataOut <= "00000000000000001110000000000000000000000000000000000000000000111000000000000000";
when "0001100010"=> dataOut <= "00000000000000000111000000000000000000000000000000000000000001110000000000000000";
when "0001100011"=> dataOut <= "00000000000000000011100000000000000000000000000000000000000011100000000000000000";
when "0001100100"=> dataOut <= "00000000000000000001110000000000000000000000000000000000000111000000000000000000";
when "0001100101"=> dataOut <= "00000000000000000000111000000000000000000000000000000000001110000000000000000000";
when "0001100110"=> dataOut <= "00000000000000000000011100000000000000000000000000000000011100000000000000000000";
when "0001100111"=> dataOut <= "00000000000000000000001110000000000000000000000000000000111000000000000000000000";
when "0001101000"=> dataOut <= "00000000000000000000000111000000000000000000000000000001110000000000000000000000";
when "0001101001"=> dataOut <= "00000000000000000000000011100000000000000000000000000011100000000000000000000000";
when "0001101010"=> dataOut <= "00000000000000000000000001110000000000000000000000000111000000000000000000000000";
when "0001101011"=> dataOut <= "00000000000000000000000000111000000000000000000000001110000000000000000000000000";
when "0001101100"=> dataOut <= "00000000000000000000000000011100000000000000000000011100000000000000000000000000";
when "0001101101"=> dataOut <= "00000000000000000000000000001110000000000000000000111000000000000000000000000000";
when "0001101110"=> dataOut <= "00000000000000000000000000000111000000000000000001110000000000000000000000000000";
when "0001101111"=> dataOut <= "00000000000000000000000000000011100000000000000011100000000000000000000000000000";
when "0001110000"=> dataOut <= "00000000000000000000000000000001110000000000000111000000000000000000000000000000";
when "0001110001"=> dataOut <= "00000000000000000000000000000000111000000000001110000000000000000000000000000000";
when "0001110010"=> dataOut <= "00000000000000000000000000000000011100000000011100000000000000000000000000000000";
when "0001110011"=> dataOut <= "00000000000000000000000000000000001110000000111000000000000000000000000000000000";
when "0001110100"=> dataOut <= "00000000000000000000000000000000000111000001110000000000000000000000000000000000";
when "0001110101"=> dataOut <= "00000000000000000000000000000000000011100011100000000000000000000000000000000000";
when "0001110110"=> dataOut <= "00000000000000000000000000000000000001110111000000000000000000000000000000000000";
when "0001110111"=> dataOut <= "00000000000000000000000000000000000000111110000000000000000000000000000000000000";
when "0001111000"=> dataOut <= "00000000000000000000000000000000000000011100000000000000000000000000000000000000";
when "0001111001"=> dataOut <= "00000000000000000000000000000000000000001000000000000000000000000000000000000000";
when "0001111010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0001111011"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";

--2
when "0010000000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0010000001"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0010000010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0010000011"=> dataOut <= "00000000000000000000000000000000000000001000000000000000000000000000000000000000";
when "0010000100"=> dataOut <= "00000000000000000000000000000000000000011100000000000000000000000000000000000000";
when "0010000101"=> dataOut <= "00000000000000000000000000000000000000111110000000000000000000000000000000000000";
when "0010000110"=> dataOut <= "00000000000000000000000000000000000001110111000000000000000000000000000000000000";
when "0010000111"=> dataOut <= "00000000000000000000000000000000000011100011100000000000000000000000000000000000";
when "0010001000"=> dataOut <= "00000000000000000000000000000000000111000001110000000000000000000000000000000000";
when "0010001001"=> dataOut <= "00000000000000000000000000000000001110001000111000000000000000000000000000000000";
when "0010001010"=> dataOut <= "00000000000000000000000000000000011100011100011100000000000000000000000000000000";
when "0010001011"=> dataOut <= "00000000000000000000000000000000111000111110001110000000000000000000000000000000";
when "0010001100"=> dataOut <= "00000000000000000000000000000001110001111111000111000000000000000000000000000000";
when "0010001101"=> dataOut <= "00000000000000000000000000000011100011111111100011100000000000000000000000000000";
when "0010001110"=> dataOut <= "00000000000000000000000000000111000111111111110001110000000000000000000000000000";
when "0010001111"=> dataOut <= "00000000000000000000000000001110001111111111111000111000000000000000000000000000";
when "0010010000"=> dataOut <= "00000000000000000000000000011100011111111111111100011100000000000000000000000000";
when "0010010001"=> dataOut <= "00000000000000000000000000111000111111111111111110001110000000000000000000000000";
when "0010010010"=> dataOut <= "00000000000000000000000001110001111111111111111111000111000000000000000000000000";
when "0010010011"=> dataOut <= "00000000000000000000000011100011111111111111111111100011100000000000000000000000";
when "0010010100"=> dataOut <= "00000000000000000000000111000111111111111111111111110001110000000000000000000000";
when "0010010101"=> dataOut <= "00000000000000000000001110001111111111111111111111111000111000000000000000000000";
when "0010010110"=> dataOut <= "00000000000000000000011100011111111111111111111111111100011100000000000000000000";
when "0010010111"=> dataOut <= "00000000000000000000111000111111111111111111111111111110001110000000000000000000";
when "0010011000"=> dataOut <= "00000000000000000001110001111111111111111111111111111111000111000000000000000000";
when "0010011001"=> dataOut <= "00000000000000000011100011111111111111111111111111111111100011100000000000000000";
when "0010011010"=> dataOut <= "00000000000000000111000111111111111111111111111111111111110001110000000000000000";
when "0010011011"=> dataOut <= "00000000000000001110001111111111111111111111111111111111111000111000000000000000";
when "0010011100"=> dataOut <= "00000000000000011100011111111111111111111111111111111111111100011100000000000000";
when "0010011101"=> dataOut <= "00000000000000111000111111111111111111111111111111111111111110001110000000000000";
when "0010011110"=> dataOut <= "00000000000001110001111111111111111111111111111111111111111111000111000000000000"; --center
when "0010011111"=> dataOut <= "00000000000000111000111111111111111111111111111111111111111110001110000000000000";
when "0010100000"=> dataOut <= "00000000000000011100011111111111111111111111111111111111111100011100000000000000";
when "0010100001"=> dataOut <= "00000000000000001110001111111111111111111111111111111111111000111000000000000000";
when "0010100010"=> dataOut <= "00000000000000000111000111111111111111111111111111111111110001110000000000000000";
when "0010100011"=> dataOut <= "00000000000000000011100011111111111111111111111111111111100011100000000000000000";
when "0010100100"=> dataOut <= "00000000000000000001110001111111111111111111111111111111000111000000000000000000";
when "0010100101"=> dataOut <= "00000000000000000000111000111111111111111111111111111110001110000000000000000000";
when "0010100110"=> dataOut <= "00000000000000000000011100011111111111111111111111111100011100000000000000000000";
when "0010100111"=> dataOut <= "00000000000000000000001110001111111111111111111111111000111000000000000000000000";
when "0010101000"=> dataOut <= "00000000000000000000000111000111111111111111111111110001110000000000000000000000";
when "0010101001"=> dataOut <= "00000000000000000000000011100011111111111111111111100011100000000000000000000000";
when "0010101010"=> dataOut <= "00000000000000000000000001110001111111111111111111000111000000000000000000000000";
when "0010101011"=> dataOut <= "00000000000000000000000000111000111111111111111110001110000000000000000000000000";
when "0010101100"=> dataOut <= "00000000000000000000000000011100011111111111111100011100000000000000000000000000";
when "0010101101"=> dataOut <= "00000000000000000000000000001110001111111111111000111000000000000000000000000000";
when "0010101110"=> dataOut <= "00000000000000000000000000000111000111111111110001110000000000000000000000000000";
when "0010101111"=> dataOut <= "00000000000000000000000000000011100011111111100011100000000000000000000000000000";
when "0010110000"=> dataOut <= "00000000000000000000000000000001110001111111000111000000000000000000000000000000";
when "0010110001"=> dataOut <= "00000000000000000000000000000000111000111110001110000000000000000000000000000000";
when "0010110010"=> dataOut <= "00000000000000000000000000000000011100011100011100000000000000000000000000000000";
when "0010110011"=> dataOut <= "00000000000000000000000000000000001110001000111000000000000000000000000000000000";
when "0010110100"=> dataOut <= "00000000000000000000000000000000000111000001110000000000000000000000000000000000";
when "0010110101"=> dataOut <= "00000000000000000000000000000000000011100011100000000000000000000000000000000000";
when "0010110110"=> dataOut <= "00000000000000000000000000000000000001110111000000000000000000000000000000000000";
when "0010110111"=> dataOut <= "00000000000000000000000000000000000000111110000000000000000000000000000000000000";
when "0010111000"=> dataOut <= "00000000000000000000000000000000000000011100000000000000000000000000000000000000";
when "0010111001"=> dataOut <= "00000000000000000000000000000000000000001000000000000000000000000000000000000000";
when "0010111010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0010111011"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";

--4
when "0100000000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0100000001"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0100000010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000111000000000000";
when "0100000011"=> dataOut <= "00000000000000000000000000000000000000001100000000000000000000000111000000000000";
when "0100000100"=> dataOut <= "00000000000000000000000000000000000000011110000000000000000000000111000000000000";
when "0100000101"=> dataOut <= "00000000000000000000000000000000000000111111000000000000000000000111000000000000";
when "0100000110"=> dataOut <= "00000000000000000000000000000000000001110011100000000000000001111111111100000000";
when "0100000111"=> dataOut <= "00000000000000000000000000000000000011100011100000000000000001111111111100000000";
when "0100001000"=> dataOut <= "00000000000000000000000000000000000111000001110000000000000001111111111100000000";
when "0100001001"=> dataOut <= "00000000000000000000000000000000001110000000111000000000000000000111000000000000";
when "0100001010"=> dataOut <= "00000000000000000000000000000000011100000000011100000000000000000111000000000000";
when "0100001011"=> dataOut <= "00000000000000000000000000000000111000000000001110000000000000000111000000000000";
when "0100001100"=> dataOut <= "00000000000000000000000000000001110000000000000111000000000000000111000000000000";
when "0100001101"=> dataOut <= "00000000000000000000000000000011100000000000000011100000000000000000000000000000";
when "0100001110"=> dataOut <= "00000000000000000000000000000111000000000000000001110000000000000000000000000000";
when "0100001111"=> dataOut <= "00000000000000000000000000001110000000000000000000111000000000000000000000000000";
when "0100010000"=> dataOut <= "00000000000000000000000000011100000000000000000000011100000000000000000000000000";
when "0100010001"=> dataOut <= "00000000000000000000000000111000000000000000000000001110000000000000000000000000";
when "0100010010"=> dataOut <= "00000000000000000000000001110000000000000000000000000111000000000000000000000000";
when "0100010011"=> dataOut <= "00000000000000000000000011100000000000000000000000000011100000000000000000000000";
when "0100010100"=> dataOut <= "00000000000000000000000111000000000000000000000000000001110000000000000000000000";
when "0100010101"=> dataOut <= "00000000000000000000001110000000000000000000000000000000111000000000000000000000";
when "0100010110"=> dataOut <= "00000000000000000000011100000000000000000000000000000000011100000000000000000000";
when "0100010111"=> dataOut <= "00000000000000000000111000000000000000000000000000000000001110000000000000000000";
when "0100011000"=> dataOut <= "00000000000000000001110000000000000000000000000000000000000111000000000000000000";
when "0100011001"=> dataOut <= "00000000000000000011100000000000000000000000000000000000000011100000000000000000";
when "0100011010"=> dataOut <= "00000000000000000111000000000000000000000000000000000000000001110000000000000000";
when "0100011011"=> dataOut <= "00000000000000001110000000000000000000000000000000000000000000111000000000000000";
when "0100011100"=> dataOut <= "00000000000000011100000000000000000000000000000000000000000000011100000000000000";
when "0100011101"=> dataOut <= "00000000000000111000000000000000000000000000000000000000000000001110000000000000";
when "0100011110"=> dataOut <= "00000000000001110000000000000000000000000000000000000000000000000111000000000000"; --center
when "0100011111"=> dataOut <= "00000000000000111000000000000000000000000000000000000000000000001110000000000000";
when "0100100000"=> dataOut <= "00000000000000011100000000000000000000000000000000000000000000011100000000000000";
when "0100100001"=> dataOut <= "00000000000000001110000000000000000000000000000000000000000000111000000000000000";
when "0100100010"=> dataOut <= "00000000000000000111000000000000000000000000000000000000000001110000000000000000";
when "0100100011"=> dataOut <= "00000000000000000011100000000000000000000000000000000000000011100000000000000000";
when "0100100100"=> dataOut <= "00000000000000000001110000000000000000000000000000000000000111000000000000000000";
when "0100100101"=> dataOut <= "00000000000000000000111000000000000000000000000000000000001110000000000000000000";
when "0100100110"=> dataOut <= "00000000000000000000011100000000000000000000000000000000011100000000000000000000";
when "0100100111"=> dataOut <= "00000000000000000000001110000000000000000000000000000000111000000000000000000000";
when "0100101000"=> dataOut <= "00000000000000000000000111000000000000000000000000000001110000000000000000000000";
when "0100101001"=> dataOut <= "00000000000000000000000011100000000000000000000000000011100000000000000000000000";
when "0100101010"=> dataOut <= "00000000000000000000000001110000000000000000000000000111000000000000000000000000";
when "0100101011"=> dataOut <= "00000000000000000000000000111000000000000000000000001110000000000000000000000000";
when "0100101100"=> dataOut <= "00000000000000000000000000011100000000000000000000011100000000000000000000000000";
when "0100101101"=> dataOut <= "00000000000000000000000000001110000000000000000000111000000000000000000000000000";
when "0100101110"=> dataOut <= "00000000000000000000000000000111000000000000000001110000000000000000000000000000";
when "0100101111"=> dataOut <= "00000000000000000000000000000011100000000000000011100000000000000000000000000000";
when "0100110000"=> dataOut <= "00000000000000000000000000000001110000000000000111000000000000000000000000000000";
when "0100110001"=> dataOut <= "00000000000000000000000000000000111000000000001110000000000000000000000000000000";
when "0100110010"=> dataOut <= "00000000000000000000000000000000011100000000011100000000000000000000000000000000";
when "0100110011"=> dataOut <= "00000000000000000000000000000000001110000000111000000000000000000000000000000000";
when "0100110100"=> dataOut <= "00000000000000000000000000000000000111000001110000000000000000000000000000000000";
when "0100110101"=> dataOut <= "00000000000000000000000000000000000011100011100000000000000000000000000000000000";
when "0100110110"=> dataOut <= "00000000000000000000000000000000000001110111000000000000000000000000000000000000";
when "0100110111"=> dataOut <= "00000000000000000000000000000000000000111110000000000000000000000000000000000000";
when "0100111000"=> dataOut <= "00000000000000000000000000000000000000011100000000000000000000000000000000000000";
when "0100111001"=> dataOut <= "00000000000000000000000000000000000000001000000000000000000000000000000000000000";
when "0100111010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0100111011"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";

--5
when "0101000000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0101000001"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0101000010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000111000000000000";
when "0101000011"=> dataOut <= "00000000000000000000000000000000000000001000000000000000000000000111000000000000";
when "0101000100"=> dataOut <= "00000000000000000000000000000000000000011100000000000000000000000111000000000000";
when "0101000101"=> dataOut <= "00000000000000000000000000000000000000111110000000000000000000000111000000000000";
when "0101000110"=> dataOut <= "00000000000000000000000000000000000001110111000000000000000001111111111100000000";
when "0101000111"=> dataOut <= "00000000000000000000000000000000000011100011100000000000000001111111111100000000";
when "0101001000"=> dataOut <= "00000000000000000000000000000000000111000001110000000000000001111111111100000000";
when "0101001001"=> dataOut <= "00000000000000000000000000000000001110001000111000000000000000000111000000000000";
when "0101001010"=> dataOut <= "00000000000000000000000000000000011100011100011100000000000000000111000000000000";
when "0101001011"=> dataOut <= "00000000000000000000000000000000111000111110001110000000000000000111000000000000";
when "0101001100"=> dataOut <= "00000000000000000000000000000001110001111111000111000000000000000111000000000000";
when "0101001101"=> dataOut <= "00000000000000000000000000000011100011111111100011100000000000000000000000000000";
when "0101001110"=> dataOut <= "00000000000000000000000000000111000111111111110001110000000000000000000000000000";
when "0101001111"=> dataOut <= "00000000000000000000000000001110001111111111111000111000000000000000000000000000";
when "0101010000"=> dataOut <= "00000000000000000000000000011100011111111111111100011100000000000000000000000000";
when "0101010001"=> dataOut <= "00000000000000000000000000111000111111111111111110001110000000000000000000000000";
when "0101010010"=> dataOut <= "00000000000000000000000001110001111111111111111111000111000000000000000000000000";
when "0101010011"=> dataOut <= "00000000000000000000000011100011111111111111111111100011100000000000000000000000";
when "0101010100"=> dataOut <= "00000000000000000000000111000111111111111111111111110001110000000000000000000000";
when "0101010101"=> dataOut <= "00000000000000000000001110001111111111111111111111111000111000000000000000000000";
when "0101010110"=> dataOut <= "00000000000000000000011100011111111111111111111111111100011100000000000000000000";
when "0101010111"=> dataOut <= "00000000000000000000111000111111111111111111111111111110001110000000000000000000";
when "0101011000"=> dataOut <= "00000000000000000001110001111111111111111111111111111111000111000000000000000000";
when "0101011001"=> dataOut <= "00000000000000000011100011111111111111111111111111111111100011100000000000000000";
when "0101011010"=> dataOut <= "00000000000000000111000111111111111111111111111111111111110001110000000000000000";
when "0101011011"=> dataOut <= "00000000000000001110001111111111111111111111111111111111111000111000000000000000";
when "0101011100"=> dataOut <= "00000000000000011100011111111111111111111111111111111111111100011100000000000000";
when "0101011101"=> dataOut <= "00000000000000111000111111111111111111111111111111111111111110001110000000000000";
when "0101011110"=> dataOut <= "00000000000001110001111111111111111111111111111111111111111111000111000000000000"; --center
when "0101011111"=> dataOut <= "00000000000000111000111111111111111111111111111111111111111110001110000000000000";
when "0101100000"=> dataOut <= "00000000000000011100011111111111111111111111111111111111111100011100000000000000";
when "0101100001"=> dataOut <= "00000000000000001110001111111111111111111111111111111111111000111000000000000000";
when "0101100010"=> dataOut <= "00000000000000000111000111111111111111111111111111111111110001110000000000000000";
when "0101100011"=> dataOut <= "00000000000000000011100011111111111111111111111111111111100011100000000000000000";
when "0101100100"=> dataOut <= "00000000000000000001110001111111111111111111111111111111000111000000000000000000";
when "0101100101"=> dataOut <= "00000000000000000000111000111111111111111111111111111110001110000000000000000000";
when "0101100110"=> dataOut <= "00000000000000000000011100011111111111111111111111111100011100000000000000000000";
when "0101100111"=> dataOut <= "00000000000000000000001110001111111111111111111111111000111000000000000000000000";
when "0101101000"=> dataOut <= "00000000000000000000000111000111111111111111111111110001110000000000000000000000";
when "0101101001"=> dataOut <= "00000000000000000000000011100011111111111111111111100011100000000000000000000000";
when "0101101010"=> dataOut <= "00000000000000000000000001110001111111111111111111000111000000000000000000000000";
when "0101101011"=> dataOut <= "00000000000000000000000000111000111111111111111110001110000000000000000000000000";
when "0101101100"=> dataOut <= "00000000000000000000000000011100011111111111111100011100000000000000000000000000";
when "0101101101"=> dataOut <= "00000000000000000000000000001110001111111111111000111000000000000000000000000000";
when "0101101110"=> dataOut <= "00000000000000000000000000000111000111111111110001110000000000000000000000000000";
when "0101101111"=> dataOut <= "00000000000000000000000000000011100011111111100011100000000000000000000000000000";
when "0101110000"=> dataOut <= "00000000000000000000000000000001110001111111000111000000000000000000000000000000";
when "0101110001"=> dataOut <= "00000000000000000000000000000000111000111110001110000000000000000000000000000000";
when "0101110010"=> dataOut <= "00000000000000000000000000000000011100011100011100000000000000000000000000000000";
when "0101110011"=> dataOut <= "00000000000000000000000000000000001110001000111000000000000000000000000000000000";
when "0101110100"=> dataOut <= "00000000000000000000000000000000000111000001110000000000000000000000000000000000";
when "0101110101"=> dataOut <= "00000000000000000000000000000000000011100011100000000000000000000000000000000000";
when "0101110110"=> dataOut <= "00000000000000000000000000000000000001110111000000000000000000000000000000000000";
when "0101110111"=> dataOut <= "00000000000000000000000000000000000000111110000000000000000000000000000000000000";
when "0101111000"=> dataOut <= "00000000000000000000000000000000000000011100000000000000000000000000000000000000";
when "0101111001"=> dataOut <= "00000000000000000000000000000000000000001000000000000000000000000000000000000000";
when "0101111010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0101111011"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";

--8
when "1000000000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "1000000001"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "1000000010"=> dataOut <= "00000000111000000011100000000000000000000000000000000000000000000000000000000000";
when "1000000011"=> dataOut <= "00000000011100000111000000000000000000001000000000000000000000000000000000000000";
when "1000000100"=> dataOut <= "00000000001110001110000000000000000000011100000000000000000000000000000000000000";
when "1000000101"=> dataOut <= "00000000000111011100000000000000000000111110000000000000000000000000000000000000";
when "1000000110"=> dataOut <= "00000000000011111000000000000000000001110111000000000000000000000000000000000000";
when "1000000111"=> dataOut <= "00000000000001110000000000000000000011100011100000000000000000000000000000000000";
when "1000001000"=> dataOut <= "00000000000011111000000000000000000111000001110000000000000000000000000000000000";
when "1000001001"=> dataOut <= "00000000000111011100000000000000001110001000111000000000000000000000000000000000";
when "1000001010"=> dataOut <= "00000000001110001110000000000000011100011100011100000000000000000000000000000000";
when "1000001011"=> dataOut <= "00000000011100000111000000000000111000111110001110000000000000000000000000000000";
when "1000001100"=> dataOut <= "00000000111000000011100000000001110001111111000111000000000000000000000000000000";
when "1000001101"=> dataOut <= "00000000000000000000000000000011100011111111100011100000000000000000000000000000";
when "1000001110"=> dataOut <= "00000000000000000000000000000111000111111111110001110000000000000000000000000000";
when "1000001111"=> dataOut <= "00000000000000000000000000001110001111111111111000111000000000000000000000000000";
when "1000010000"=> dataOut <= "00000000000000000000000000011100011111111111111100011100000000000000000000000000";
when "1000010001"=> dataOut <= "00000000000000000000000000111000111111111111111110001110000000000000000000000000";
when "1000010010"=> dataOut <= "00000000000000000000000001110001111111111111111111000111000000000000000000000000";
when "1000010011"=> dataOut <= "00000000000000000000000011100011111111111111111111100011100000000000000000000000";
when "1000010100"=> dataOut <= "00000000000000000000000111000111111111111111111111110001110000000000000000000000";
when "1000010101"=> dataOut <= "00000000000000000000001110001111111111111111111111111000111000000000000000000000";
when "1000010110"=> dataOut <= "00000000000000000000011100011111111111111111111111111100011100000000000000000000";
when "1000010111"=> dataOut <= "00000000000000000000111000111111111111111111111111111110001110000000000000000000";
when "1000011000"=> dataOut <= "00000000000000000001110001111111111111111111111111111111000111000000000000000000";
when "1000011001"=> dataOut <= "00000000000000000011100011111111111111111111111111111111100011100000000000000000";
when "1000011010"=> dataOut <= "00000000000000000111000111111111111111111111111111111111110001110000000000000000";
when "1000011011"=> dataOut <= "00000000000000001110001111111111111111111111111111111111111000111000000000000000";
when "1000011100"=> dataOut <= "00000000000000011100011111111111111111111111111111111111111100011100000000000000";
when "1000011101"=> dataOut <= "00000000000000111000111111111111111111111111111111111111111110001110000000000000";
when "1000011110"=> dataOut <= "00000000000001110001111111111111111111111111111111111111111111000111000000000000"; --center
when "1000011111"=> dataOut <= "00000000000000111000111111111111111111111111111111111111111110001110000000000000";
when "1000100000"=> dataOut <= "00000000000000011100011111111111111111111111111111111111111100011100000000000000";
when "1000100001"=> dataOut <= "00000000000000001110001111111111111111111111111111111111111000111000000000000000";
when "1000100010"=> dataOut <= "00000000000000000111000111111111111111111111111111111111110001110000000000000000";
when "1000100011"=> dataOut <= "00000000000000000011100011111111111111111111111111111111100011100000000000000000";
when "1000100100"=> dataOut <= "00000000000000000001110001111111111111111111111111111111000111000000000000000000";
when "1000100101"=> dataOut <= "00000000000000000000111000111111111111111111111111111110001110000000000000000000";
when "1000100110"=> dataOut <= "00000000000000000000011100011111111111111111111111111100011100000000000000000000";
when "1000100111"=> dataOut <= "00000000000000000000001110001111111111111111111111111000111000000000000000000000";
when "1000101000"=> dataOut <= "00000000000000000000000111000111111111111111111111110001110000000000000000000000";
when "1000101001"=> dataOut <= "00000000000000000000000011100011111111111111111111100011100000000000000000000000";
when "1000101010"=> dataOut <= "00000000000000000000000001110001111111111111111111000111000000000000000000000000";
when "1000101011"=> dataOut <= "00000000000000000000000000111000111111111111111110001110000000000000000000000000";
when "1000101100"=> dataOut <= "00000000000000000000000000011100011111111111111100011100000000000000000000000000";
when "1000101101"=> dataOut <= "00000000000000000000000000001110001111111111111000111000000000000000000000000000";
when "1000101110"=> dataOut <= "00000000000000000000000000000111000111111111110001110000000000000000000000000000";
when "1000101111"=> dataOut <= "00000000000000000000000000000011100011111111100011100000000000000000000000000000";
when "1000110000"=> dataOut <= "00000000000000000000000000000001110001111111000111000000000000000000000000000000";
when "1000110001"=> dataOut <= "00000000000000000000000000000000111000111110001110000000000000000000000000000000";
when "1000110010"=> dataOut <= "00000000000000000000000000000000011100011100011100000000000000000000000000000000";
when "1000110011"=> dataOut <= "00000000000000000000000000000000001110001000111000000000000000000000000000000000";
when "1000110100"=> dataOut <= "00000000000000000000000000000000000111000001110000000000000000000000000000000000";
when "1000110101"=> dataOut <= "00000000000000000000000000000000000011100011100000000000000000000000000000000000";
when "1000110110"=> dataOut <= "00000000000000000000000000000000000001110111000000000000000000000000000000000000";
when "1000110111"=> dataOut <= "00000000000000000000000000000000000000111110000000000000000000000000000000000000";
when "1000111000"=> dataOut <= "00000000000000000000000000000000000000011100000000000000000000000000000000000000";
when "1000111001"=> dataOut <= "00000000000000000000000000000000000000001000000000000000000000000000000000000000";
when "1000111010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "1000111011"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";

--11
when "1011000000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "1011000001"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "1011000010"=> dataOut <= "00000000111000000011100000000000000000000000000000000000000000000111000000000000";
when "1011000011"=> dataOut <= "00000000011100000111000000000000000000001000000000000000000000000111000000000000";
when "1011000100"=> dataOut <= "00000000001110001110000000000000000000011100000000000000000000000111000000000000";
when "1011000101"=> dataOut <= "00000000000111011100000000000000000000111110000000000000000000000111000000000000";
when "1011000110"=> dataOut <= "00000000000011111000000000000000000001110111000000000000000000111111111000000000";
when "1011000111"=> dataOut <= "00000000000001110000000000000000000011100011100000000000000000111111111000000000";
when "1011001000"=> dataOut <= "00000000000011111000000000000000000111000001110000000000000000111111111000000000";
when "1011001001"=> dataOut <= "00000000000111011100000000000000001110001000111000000000000000000111000000000000";
when "1011001010"=> dataOut <= "00000000001110001110000000000000011100011100011100000000000000000111000000000000";
when "1011001011"=> dataOut <= "00000000011100000111000000000000111000111110001110000000000000000111000000000000";
when "1011001100"=> dataOut <= "00000000111000000011100000000001110001111111000111000000000000000111000000000000";
when "1011001101"=> dataOut <= "00000000000000000000000000000011100011111111100011100000000000000000000000000000";
when "1011001110"=> dataOut <= "00000000000000000000000000000111000111111111110001110000000000000000000000000000";
when "1011001111"=> dataOut <= "00000000000000000000000000001110001111111111111000111000000000000000000000000000";
when "1011010000"=> dataOut <= "00000000000000000000000000011100011111111111111100011100000000000000000000000000";
when "1011010001"=> dataOut <= "00000000000000000000000000111000111111111111111110001110000000000000000000000000";
when "1011010010"=> dataOut <= "00000000000000000000000001110001111111111111111111000111000000000000000000000000";
when "1011010011"=> dataOut <= "00000000000000000000000011100011111111111111111111100011100000000000000000000000";
when "1011010100"=> dataOut <= "00000000000000000000000111000111111111111111111111110001110000000000000000000000";
when "1011010101"=> dataOut <= "00000000000000000000001110001111111111111111111111111000111000000000000000000000";
when "1011010110"=> dataOut <= "00000000000000000000011100011111111111111111111111111100011100000000000000000000";
when "1011010111"=> dataOut <= "00000000000000000000111000111111111111111111111111111110001110000000000000000000";
when "1011011000"=> dataOut <= "00000000000000000001110001111111111111111111111111111111000111000000000000000000";
when "1011011001"=> dataOut <= "00000000000000000011100011111111111111111111111111111111100011100000000000000000";
when "1011011010"=> dataOut <= "00000000000000000111000111111111111111111111111111111111110001110000000000000000";
when "1011011011"=> dataOut <= "00000000000000001110001111111111111111111111111111111111111000111000000000000000";
when "1011011100"=> dataOut <= "00000000000000011100011111111111111111111111111111111111111100011100000000000000";
when "1011011101"=> dataOut <= "00000000000000111000111111111111111111111111111111111111111110001110000000000000";
when "1011011110"=> dataOut <= "00000000000001110001111111111111111111111111111111111111111111000111000000000000"; --center
when "1011011111"=> dataOut <= "00000000000000111000111111111111111111111111111111111111111110001110000000000000";
when "1011100000"=> dataOut <= "00000000000000011100011111111111111111111111111111111111111100011100000000000000";
when "1011100001"=> dataOut <= "00000000000000001110001111111111111111111111111111111111111000111000000000000000";
when "1011100010"=> dataOut <= "00000000000000000111000111111111111111111111111111111111110001110000000000000000";
when "1011100011"=> dataOut <= "00000000000000000011100011111111111111111111111111111111100011100000000000000000";
when "1011100100"=> dataOut <= "00000000000000000001110001111111111111111111111111111111000111000000000000000000";
when "1011100101"=> dataOut <= "00000000000000000000111000111111111111111111111111111110001110000000000000000000";
when "1011100110"=> dataOut <= "00000000000000000000011100011111111111111111111111111100011100000000000000000000";
when "1011100111"=> dataOut <= "00000000000000000000001110001111111111111111111111111000111000000000000000000000";
when "1011101000"=> dataOut <= "00000000000000000000000111000111111111111111111111110001110000000000000000000000";
when "1011101001"=> dataOut <= "00000000000000000000000011100011111111111111111111100011100000000000000000000000";
when "1011101010"=> dataOut <= "00000000000000000000000001110001111111111111111111000111000000000000000000000000";
when "1011101011"=> dataOut <= "00000000000000000000000000111000111111111111111110001110000000000000000000000000";
when "1011101100"=> dataOut <= "00000000000000000000000000011100011111111111111100011100000000000000000000000000";
when "1011101101"=> dataOut <= "00000000000000000000000000001110001111111111111000111000000000000000000000000000";
when "1011101110"=> dataOut <= "00000000000000000000000000000111000111111111110001110000000000000000000000000000";
when "1011101111"=> dataOut <= "00000000000000000000000000000011100011111111100011100000000000000000000000000000";
when "1011110000"=> dataOut <= "00000000000000000000000000000001110001111111000111000000000000000000000000000000";
when "1011110001"=> dataOut <= "00000000000000000000000000000000111000111110001110000000000000000000000000000000";
when "1011110010"=> dataOut <= "00000000000000000000000000000000011100011100011100000000000000000000000000000000";
when "1011110011"=> dataOut <= "00000000000000000000000000000000001110001000111000000000000000000000000000000000";
when "1011110100"=> dataOut <= "00000000000000000000000000000000000111000001110000000000000000000000000000000000";
when "1011110101"=> dataOut <= "00000000000000000000000000000000000011100011100000000000000000000000000000000000";
when "1011110110"=> dataOut <= "00000000000000000000000000000000000001110111000000000000000000000000000000000000";
when "1011110111"=> dataOut <= "00000000000000000000000000000000000000111110000000000000000000000000000000000000";
when "1011111000"=> dataOut <= "00000000000000000000000000000000000000011100000000000000000000000000000000000000";
when "1011111001"=> dataOut <= "00000000000000000000000000000000000000001000000000000000000000000000000000000000";
when "1011111010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "1011111011"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";

when others => dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
end case;
end process;
end RTL;