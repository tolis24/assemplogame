library ieee;
use ieee.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity icon_rom is
port (countV : in std_logic_vector(9 downto 0);
		pointer : in std_logic_vector(3 downto 0);
		dataOut : out std_logic_vector(79 downto 0));
end icon_rom;

architecture RTL of icon_rom is

signal row : std_logic_vector(9 downto 0);
signal address : std_logic_vector(9 downto 0);

begin

process (countV)
begin 
	if unsigned(countV) < 60 then 
		row <= countV;
	elsif unsigned(countV) < 120 then
		row <= unsigned(countV) - 60;
	elsif unsigned(countV) < 180 then
		row <= unsigned(countV) - 120;
	elsif unsigned(countV) < 240 then
		row <= unsigned(countV) - 180;
	elsif unsigned(countV) < 300 then
		row <= unsigned(countV) - 240;
	elsif unsigned(countV) < 360 then
		row <= unsigned(countV) - 300;
	elsif unsigned(countV) < 420 then
		row <= unsigned(countV) - 360;
	elsif unsigned(countV) < 480 then
		row <= unsigned(countV) - 420;
	else
		row <= (others => '0');
	end if;
end process;

		
address(9 downto 6) <= pointer;
address(5 downto 0) <= row(5 downto 0);

process(address)
begin
case address is
-- 0
when "0000000000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000000001"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000000010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000000011"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000000100"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000000101"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000000110"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000000111"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000001000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000001001"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000001010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000001011"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000001100"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000001101"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000001110"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000001111"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000010000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000010001"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000010010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000010011"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000010100"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000010101"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000010110"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000010111"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000011000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000011001"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000011010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000011011"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000011100"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000011101"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000011110"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000011111"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000100000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000100001"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000100010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000100011"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000100100"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000100101"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000100110"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000100111"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000101000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000101001"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000101010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000101011"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000101100"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000101101"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000101110"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000101111"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000110000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000110001"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000110010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000110011"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000110100"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000110101"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000110110"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000110111"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000111000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000111001"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";
when "0000111010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0000111011"=> dataOut <= "11111111111111111111111111111111111111111111111111111111111111111111111111111111";

--1
when "0001000000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0001000001"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0001000010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0001000011"=> dataOut <= "00000000000000000000000000000000000000001000000000000000000000000000000000000000";
when "0001000100"=> dataOut <= "00000000000000000000000000000000000000011100000000000000000000000000000000000000";
when "0001000101"=> dataOut <= "00000000000000000000000000000000000000111110000000000000000000000000000000000000";
when "0001000110"=> dataOut <= "00000000000000000000000000000000000001110111000000000000000000000000000000000000";
when "0001000111"=> dataOut <= "00000000000000000000000000000000000011100111000000000000000000000000000000000000";
when "0001001000"=> dataOut <= "00000000000000000000000000000000000111000011100000000000000000000000000000000000";
when "0001001001"=> dataOut <= "00000000000000000000000000000000001110000001110000000000000000000000000000000000";
when "0001001010"=> dataOut <= "00000000000000000000000000000000011100000000111000000000000000000000000000000000";
when "0001001011"=> dataOut <= "00000000000000000000000000000000111000000000011100000000000000000000000000000000";
when "0001001100"=> dataOut <= "00000000000000000000000000000001110000000000001110000000000000000000000000000000";
when "0001001101"=> dataOut <= "00000000000000000000000000000011100000000000000111000000000000000000000000000000";
when "0001001110"=> dataOut <= "00000000000000000000000000000111000000000000000011100000000000000000000000000000";
when "0001001111"=> dataOut <= "00000000000000000000000000001110000000000000000001110000000000000000000000000000";
when "0001010000"=> dataOut <= "00000000000000000000000000011100000000000000000000111000000000000000000000000000";
when "0001010001"=> dataOut <= "00000000000000000000000000111000000000000000000000011100000000000000000000000000";
when "0001010010"=> dataOut <= "00000000000000000000000001110000000000000000000000001110000000000000000000000000";
when "0001010011"=> dataOut <= "00000000000000000000000011100000000000000000000000000111000000000000000000000000";
when "0001010100"=> dataOut <= "00000000000000000000000111000000000000000000000000000011100000000000000000000000";
when "0001010101"=> dataOut <= "00000000000000000000001110000000000000000000000000000001110000000000000000000000";
when "0001010110"=> dataOut <= "00000000000000000000011100000000000000000000000000000000111000000000000000000000";
when "0001010111"=> dataOut <= "00000000000000000000111000000000000000000000000000000000011100000000000000000000";
when "0001011000"=> dataOut <= "00000000000000000001110000000000000000000000000000000000001110000000000000000000";
when "0001011001"=> dataOut <= "00000000000000000011100000000000000000000000000000000000000111000000000000000000";
when "0001011010"=> dataOut <= "00000000000000000111000000000000000000000000000000000000000011100000000000000000";
when "0001011011"=> dataOut <= "00000000000000001110000000000000000000000000000000000000000001110000000000000000";
when "0001011100"=> dataOut <= "00000000000000011100000000000000000000000000000000000000000000111000000000000000";
when "0001011101"=> dataOut <= "00000000000000111000000000000000000000000000000000000000000000011100000000000000";
when "0001011110"=> dataOut <= "00000000000001110000000000000000000000000000000000000000000000001110000000000000"; --center
when "0001011111"=> dataOut <= "00000000000000111000000000000000000000000000000000000000000000011100000000000000";
when "0001100000"=> dataOut <= "00000000000000011100000000000000000000000000000000000000000000111000000000000000";
when "0001100001"=> dataOut <= "00000000000000001110000000000000000000000000000000000000000001110000000000000000";
when "0001100010"=> dataOut <= "00000000000000000111000000000000000000000000000000000000000011100000000000000000";
when "0001100011"=> dataOut <= "00000000000000000011100000000000000000000000000000000000000111000000000000000000";
when "0001100100"=> dataOut <= "00000000000000000001110000000000000000000000000000000000001110000000000000000000";
when "0001100101"=> dataOut <= "00000000000000000000111000000000000000000000000000000000011100000000000000000000";
when "0001100110"=> dataOut <= "00000000000000000000011100000000000000000000000000000000111000000000000000000000";
when "0001100111"=> dataOut <= "00000000000000000000001110000000000000000000000000000001110000000000000000000000";
when "0001101000"=> dataOut <= "00000000000000000000000111000000000000000000000000000011100000000000000000000000";
when "0001101001"=> dataOut <= "00000000000000000000000011100000000000000000000000000111000000000000000000000000";
when "0001101010"=> dataOut <= "00000000000000000000000001110000000000000000000000001110000000000000000000000000";
when "0001101011"=> dataOut <= "00000000000000000000000000111000000000000000000000011100000000000000000000000000";
when "0001101100"=> dataOut <= "00000000000000000000000000011100000000000000000000111000000000000000000000000000";
when "0001101101"=> dataOut <= "00000000000000000000000000001110000000000000000001110000000000000000000000000000";
when "0001101110"=> dataOut <= "00000000000000000000000000000111000000000000000011100000000000000000000000000000";
when "0001101111"=> dataOut <= "00000000000000000000000000000011100000000000000111000000000000000000000000000000";
when "0001110000"=> dataOut <= "00000000000000000000000000000001110000000000001110000000000000000000000000000000";
when "0001110001"=> dataOut <= "00000000000000000000000000000000111000000000011100000000000000000000000000000000";
when "0001110010"=> dataOut <= "00000000000000000000000000000000011100000000111000000000000000000000000000000000";
when "0001110011"=> dataOut <= "00000000000000000000000000000000001110000001110000000000000000000000000000000000";
when "0001110100"=> dataOut <= "00000000000000000000000000000000000111000011100000000000000000000000000000000000";
when "0001110101"=> dataOut <= "00000000000000000000000000000000000011100111000000000000000000000000000000000000";
when "0001110110"=> dataOut <= "00000000000000000000000000000000000001110111000000000000000000000000000000000000";
when "0001110111"=> dataOut <= "00000000000000000000000000000000000000111110000000000000000000000000000000000000";
when "0001111000"=> dataOut <= "00000000000000000000000000000000000000011100000000000000000000000000000000000000";
when "0001111001"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0001111010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0001111011"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";

--2
when "0010000000"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0010000001"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0010000010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0010000011"=> dataOut <= "00000000000000000000000000000000000000001000000000000000000000000000000000000000";
when "0010000100"=> dataOut <= "00000000000000000000000000000000000000011100000000000000000000000000000000000000";
when "0010000101"=> dataOut <= "00000000000000000000000000000000000000111110000000000000000000000000000000000000";
when "0010000110"=> dataOut <= "00000000000000000000000000000000000001110111000000000000000000000000000000000000";
when "0010000111"=> dataOut <= "00000000000000000000000000000000000011100111000000000000000000000000000000000000";
when "0010001000"=> dataOut <= "00000000000000000000000000000000000111000011100000000000000000000000000000000000";
when "0010001001"=> dataOut <= "00000000000000000000000000000000001110001001110000000000000000000000000000000000";
when "0010001010"=> dataOut <= "00000000000000000000000000000000011100001000111000000000000000000000000000000000";
when "0010001011"=> dataOut <= "00000000000000000000000000000000111000011100011100000000000000000000000000000000";
when "0010001100"=> dataOut <= "00000000000000000000000000000001110001111110001110000000000000000000000000000000";
when "0010001101"=> dataOut <= "00000000000000000000000000000011100011111111000111000000000000000000000000000000";
when "0010001110"=> dataOut <= "00000000000000000000000000000111000111111111100011100000000000000000000000000000";
when "0010001111"=> dataOut <= "00000000000000000000000000001110000111111111110001110000000000000000000000000000";
when "0010010000"=> dataOut <= "00000000000000000000000000011100011111111111111000111000000000000000000000000000";
when "0010010001"=> dataOut <= "00000000000000000000000000111000111111111111111100011100000000000000000000000000";
when "0010010010"=> dataOut <= "00000000000000000000000001110001111111111111111110001110000000000000000000000000";
when "0010010011"=> dataOut <= "00000000000000000000000011100011111111111111111111000111000000000000000000000000";
when "0010010100"=> dataOut <= "00000000000000000000000111000111111111111111111111100011100000000000000000000000";
when "0010010101"=> dataOut <= "00000000000000000000001110001111111111111111111111110001110000000000000000000000";
when "0010010110"=> dataOut <= "00000000000000000000011100011111111111111111111111111000111000000000000000000000";
when "0010010111"=> dataOut <= "00000000000000000000111000111111111111111111111111111100011100000000000000000000";
when "0010011000"=> dataOut <= "00000000000000000001110001111111111111111111111111111110001110000000000000000000";
when "0010011001"=> dataOut <= "00000000000000000011100011111111111111111111111111111111000111000000000000000000";
when "0010011010"=> dataOut <= "00000000000000000111000111111111111111111111111111111111100011100000000000000000";
when "0010011011"=> dataOut <= "00000000000000001110001111111111111111111111111111111111110001110000000000000000";
when "0010011100"=> dataOut <= "00000000000000011100011111111111111111111111111111111111111000111000000000000000";
when "0010011101"=> dataOut <= "00000000000000111000111111111111111111111111111111111111111100011100000000000000";
when "0010011110"=> dataOut <= "00000000000001110001111111111111111111111111111111111111111110001110000000000000"; --center
when "0010011111"=> dataOut <= "00000000000000111000111111111111111111111111111111111111111100011100000000000000";
when "0010100000"=> dataOut <= "00000000000000011100011111111111111111111111111111111111111000111000000000000000";
when "0010100001"=> dataOut <= "00000000000000001110001111111111111111111111111111111111110001110000000000000000";
when "0010100010"=> dataOut <= "00000000000000000111000111111111111111111111111111111111100011100000000000000000";
when "0010100011"=> dataOut <= "00000000000000000011100011111111111111111111111111111111000111000000000000000000";
when "0010100100"=> dataOut <= "00000000000000000001110001111111111111111111111111111110001110000000000000000000";
when "0010100101"=> dataOut <= "00000000000000000000111000111111111111111111111111111100011100000000000000000000";
when "0010100110"=> dataOut <= "00000000000000000000011100011111111111111111111111111000111000000000000000000000";
when "0010100111"=> dataOut <= "00000000000000000000001110001111111111111111111111110001110000000000000000000000";
when "0010101000"=> dataOut <= "00000000000000000000000111000111111111111111111111100011100000000000000000000000";
when "0010101001"=> dataOut <= "00000000000000000000000011100011111111111111111111000111000000000000000000000000";
when "0010101010"=> dataOut <= "00000000000000000000000001110001111111111111111110001110000000000000000000000000";
when "0010101011"=> dataOut <= "00000000000000000000000000111000111111111111111100011100000000000000000000000000";
when "0010101100"=> dataOut <= "00000000000000000000000000011100011111111111111000111000000000000000000000000000";
when "0010101101"=> dataOut <= "00000000000000000000000000001110001111111111110001110000000000000000000000000000";
when "0010101110"=> dataOut <= "00000000000000000000000000000111000111111111100011100000000000000000000000000000";
when "0010101111"=> dataOut <= "00000000000000000000000000000011100011111111000111000000000000000000000000000000";
when "0010110000"=> dataOut <= "00000000000000000000000000000001110001111110001110000000000000000000000000000000";
when "0010110001"=> dataOut <= "00000000000000000000000000000000111000111100011100000000000000000000000000000000";
when "0010110010"=> dataOut <= "00000000000000000000000000000000011100011000111000000000000000000000000000000000";
when "0010110011"=> dataOut <= "00000000000000000000000000000000001110001001110000000000000000000000000000000000";
when "0010110100"=> dataOut <= "00000000000000000000000000000000000111000011100000000000000000000000000000000000";
when "0010110101"=> dataOut <= "00000000000000000000000000000000000011100111000000000000000000000000000000000000";
when "0010110110"=> dataOut <= "00000000000000000000000000000000000001110111000000000000000000000000000000000000";
when "0010110111"=> dataOut <= "00000000000000000000000000000000000000111110000000000000000000000000000000000000";
when "0010111000"=> dataOut <= "00000000000000000000000000000000000000011100000000000000000000000000000000000000";
when "0010111001"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0010111010"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
when "0010111011"=> dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";


when others => dataOut <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
end case;
end process;
end RTL;